// Note the Verilog-1995 module declaration syntax here:
module top_module(clk, reset, in, out);
    input clk;
    input reset;    // Synchronous reset to state B
    input in;
    output out;//  
    reg out;

    reg present_state, next_state;
    parameter A= 0, B=1;

    always @(posedge clk) begin
        if (reset) begin  
            present_state <= B;
        end else 
            begin
                 present_state <= next_state; 
            end
    end
    
    always@(*) begin
            case (present_state)
                // Fill in state transition logic
                A: next_state = in? A: B;
                B: next_state = in? B: A;   
            endcase
    end

    assign out = (present_state == A)? 0:1;
endmodule
